//-----------------------------------------------------------
// Author        : Jzhen
// Email         : majx1996@outlook.com
// Last modified : 2023-04-24 00:42
// Filename      : axi_si.v
// Description   : 
//-----------------------------------------------------------
module axi_si();

























endmodule
